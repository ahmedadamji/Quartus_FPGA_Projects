module SimpleLogic  (
	A,
	B,
	Out
);

	input A;
	input B;
	
	output Out;
	
	and(Out, A, B);
	



endmodule