module OrGate  (
	A,
	B,
	Out
);

	input A;
	input B;
	
	output Out;
	
	or(Out, A, B);
	



endmodule 